library ieee;
use ieee.std_logic_1164.all;

entity Mux2_1minutos is
port( Sel: in std_logic;
		D0, D1: in std_logic_vector (5 downto 0);
		Q: out std_logic_vector (5 downto 0));
end Mux2_1minutos;

architecture desarrollo of Mux2_1minutos is
signal temp: std_logic_vector (5 downto 0);
begin
	process(Sel)
	begin
		case Sel is
			when '0' => temp<=D0;
			when '1' => temp<=D1;
		end case;
	end process;
Q<=temp;
end desarrollo;